// rename/dispatch shit
module dispatcher
    import rv32i_types::*;
    #(
        parameter SS = 2,
        parameter PR_ENTRIES = 64,
        parameter ROB_DEPTH = 8
    )
    (
        input logic clk, 
        input logic rst,

        // inform inst queue to pop another inst 
        output logic pop_inst_q, 
        output logic avail_inst, 
        // This is based on whether the reservation station is full or not
        input logic alu_table_full, 
        input logic mult_table_full, 
        input instruction_info_reg_t view_inst_tail [SS], 
        input logic inst_q_empty, 
        input logic rob_full,

        // inst input from the inst queue
        input instruction_info_reg_t inst [SS],

        // Acquire RAT Mapping
        output logic [4:0] isa_rs1 [SS], 
        output logic [4:0] isa_rs2 [SS], 
        // Width of the phys. reg. is larger because we're supporting twice 
        // as many internal phys. reg as arch. reg. 
        input logic [5:0] rat_rs1 [SS], 
        input logic [5:0] rat_rs2 [SS], 

        // Phys Reg to Update Mapping for
        output logic [4:0] isa_rd[SS],
        // New Phys RD for ISA RD
        output logic [5:0] rat_rd[SS],

        // Acquire new mapping for destination register 
        // Free list is popped same time that the inst queue is popped
        input logic [5:0] free_rat_rds [SS], 

        // Physical register ports 
        output physical_reg_request_t dispatch_request [SS],
        input physical_reg_response_t dispatch_reg_data [SS],

        // Acquire ROB_ID for current inst. 
        // This will be useful for updating the reservation station later
        input logic [$clog2(ROB_DEPTH)-1:0] rob_id_next [SS],
        
        // Build a super dispatch struct to feed into the ROB and the Reservation Station
        output super_dispatch_t rs_rob_entry [SS],
        output logic [1:0] update_rat, 

        input logic lsq_full
    ); 

    // We want to gain new input every clock cycle from the free list and inst queues
    // unless we need to stall because of backlog in the reservation station 
    // Because this signal will drive popping from two queues, ensure that if the inst. queue is 
    // empty, then we don't still pop from the free list queue
    // We latch this signal because we want this signal to be 0 when rst is high
    always_ff @ (posedge clk) begin
        if(rst) begin
            avail_inst <= '0; 
        end
        else begin
            avail_inst <= pop_inst_q; 
        end
    end

    // assign update_rat = avail_inst && inst[0].has_rd;
    // if both the tables are available OR if the multiplication table is not available but the next two insructions are addition based
    assign pop_inst_q = ~inst_q_empty && ~rob_full && ~lsq_full && 
    ((~alu_table_full && ~mult_table_full) || (alu_table_full && (view_inst_tail[0].is_mul && view_inst_tail[1].is_mul)) || (mult_table_full && (~view_inst_tail[0].is_mul && ~view_inst_tail[1].is_mul))); 
    logic alpha; 
    assign alpha = ~inst_q_empty && ~rob_full && ~(alu_table_full || mult_table_full);
    
    always_comb begin
        if(avail_inst) begin
            // need to build rat signals, rvfi signals
            // if the second way source registers depend on the first way destination registers, the CDB will directly update those
            // if the first way source registers depend on the last pair's second way's destination register the mappings should be intact
            // if two instructions in the same way write to the same isa, then the first way shouldn't update the rat
            // if two instructions, one in the second way of the previous pair, then both should update the rat 

            for(int i = 0; i < SS; i++) begin
                if(avail_inst && inst[i].has_rd && (inst[i].rd_s != '0)) begin
                    // if two instructions in the same way write to the same isa, then the first way shouldn't update the rat
                    update_rat[i] = '1; 
                    if((i == 0) && (isa_rd[1] == isa_rd[0])) begin
                        update_rat[i] = '0; 
                    end
                end
                else begin
                    update_rat[i] = '0; 
                end
                // Get the ISA Regs to read
                isa_rs1[i] = inst[i].rs1_s;
                isa_rs2[i] = inst[i].rs2_s;
                // Set the RAT Entry whose mapping to update with free list
                isa_rd[i] = inst[i].rd_s;
                rat_rd[i] = free_rat_rds[i];
                // Set the inputs to the phys. reg. file that we would like to read
                // We get the phys. eg. to read from by the RAT
                // dispatch_request[i].rs1_s = rat_rs1[i];
                // dispatch_request[i].rs2_s = rat_rs2[i];
                if(inst[i].has_rd && inst[i].rd_s != '0) begin
                    dispatch_request[i].rd_s = free_rat_rds[i];
                    dispatch_request[i].rd_en = 1'b1;
                end
                else begin
                    dispatch_request[i].rd_s = '0;
                    dispatch_request[i].rd_en = 1'b0;
                end
                dispatch_request[i].rd_v.register_value = 'x;
                dispatch_request[i].rd_v.ROB_ID = rob_id_next[i];
                dispatch_request[i].rd_v.dependency = 'x;


                // ROB Setup
                rs_rob_entry[i].rob.rob_id = rob_id_next[i];
                rs_rob_entry[i].rob.commit = 1'b0;
                rs_rob_entry[i].rob.branch_enable = 'x;
                rs_rob_entry[i].rob.mispredict = '0;
                rs_rob_entry[i].rs_entry.rs1_source = dispatch_reg_data[i].rs1_v.ROB_ID;
                rs_rob_entry[i].rs_entry.rs2_source = dispatch_reg_data[i].rs2_v.ROB_ID;
                rs_rob_entry[i].rs_entry.full = 1'b0; // Mark as effectively empty

                
                if(i == 1 && (isa_rs1[1] == isa_rd[0]) && (isa_rs1[1] != '0)) begin
                    dispatch_request[i].rs1_s = rat_rd[0];
                    rs_rob_entry[i].rat.rs1 = rat_rd[0]; 
                    rs_rob_entry[i].rs_entry.rs1_source = rob_id_next[0];
                end
                else begin
                    rs_rob_entry[i].rat.rs1 = rat_rs1[i];
                    dispatch_request[i].rs1_s = rat_rs1[i];
                end
                if(i == 1 && (isa_rs2[1] == isa_rd[0]) && (isa_rs2[1] != '0)) begin
                    dispatch_request[i].rs2_s = rat_rd[0]; 
                    rs_rob_entry[i].rat.rs2 = rat_rd[0]; 
                    rs_rob_entry[i].rs_entry.rs2_source = rob_id_next[0];
                end
                else begin
                    dispatch_request[i].rs2_s = rat_rs2[i];
                    rs_rob_entry[i].rat.rs2 = rat_rs2[i];
                end

                if(i == 1 && (isa_rs1[1] == isa_rd[0]) && (isa_rs1[1] != '0)) begin
                    rs_rob_entry[i].rs_entry.input1_met = '0;  
                end 
                else if(~inst[i].execute_operand1[0] || inst[i].is_branch || inst[i].is_jump) begin
                    rs_rob_entry[i].rs_entry.input1_met = ~dispatch_reg_data[i].rs1_v.dependency; 
                end
                else begin
                    rs_rob_entry[i].rs_entry.input1_met = '1;  
                end

                if(i == 1 && (isa_rs2[1] == isa_rd[0]) && (isa_rs2[1] != '0)) begin
                    rs_rob_entry[i].rs_entry.input2_met = '0; 
                end
                else if(~inst[i].execute_operand2[0] || inst[i].is_branch || inst[i].is_jump) begin
                    rs_rob_entry[i].rs_entry.input2_met = ~dispatch_reg_data[i].rs2_v.dependency; 
                end
                else begin
                    rs_rob_entry[i].rs_entry.input2_met = '1; 
                end


                // RVFI Setup
                rs_rob_entry[i].rvfi.valid = inst[i].valid;
                rs_rob_entry[i].rvfi.order = 'x; // Determine order in ROB 
                rs_rob_entry[i].rvfi.inst = inst[i].inst;
                rs_rob_entry[i].rvfi.rs1_addr = inst[i].rs1_s;
                rs_rob_entry[i].rvfi.rs2_addr = inst[i].rs2_s;
                rs_rob_entry[i].rvfi.rs1_rdata = 'x;
                rs_rob_entry[i].rvfi.rs2_rdata = 'x;
                rs_rob_entry[i].rvfi.rd_addr = inst[i].rd_s;
                rs_rob_entry[i].rvfi.rd_wdata = 'x;
                rs_rob_entry[i].rvfi.pc_rdata = inst[i].pc_curr;
                rs_rob_entry[i].rvfi.pc_wdata = inst[i].pc_next;
                rs_rob_entry[i].rvfi.mem_addr = 'x;
                // Need to compute rmask/wmask based on type of mem op
                // By default we don't make a memory request
                rs_rob_entry[i].rvfi.mem_rmask = inst[i].rmask;
                rs_rob_entry[i].rvfi.mem_wmask = inst[i].wmask;
                rs_rob_entry[i].rvfi.mem_rdata = 'x;
                rs_rob_entry[i].rvfi.mem_wdata = 'x;
                
                //inst setup
                rs_rob_entry[i].inst = inst[i];

                //Rat Registers
                // If ISA is R0, then since we don't update the RAT we'll always get rat_r = PR0
                // The only issue is we pop a free list reg regardless which could cause problems
                // rs_rob_entry[i].rat.rs1 = rat_rs1[i];
                // rs_rob_entry[i].rat.rs2 = rat_rs2[i];
                // Don't need to save the mapping we are overwritting because that is in the RRAT
                if(inst[i].has_rd && inst[i].rd_s != '0)
                    rs_rob_entry[i].rat.rd = free_rat_rds[i];
                else
                    rs_rob_entry[i].rat.rd = '0;

                // Set cross tail for load store queue
                rs_rob_entry[i].cross_entry = 'x;
            end
        end
        else begin
            for(int i = 0; i < SS; i++) begin
                update_rat[i] = '0; 
                isa_rs1[i] = 'x;
                isa_rs2[i] = 'x;
                isa_rd[i] = 'x;
                rat_rd[i] = 'x;
                // Set the inputs to the phys. reg. file that we would like to read
                // We get the phys. eg. to read from by the RAT
                dispatch_request[i].rs1_s = 'x; 
                dispatch_request[i].rs2_s = 'x;
                dispatch_request[i].rd_s = 'x;
                dispatch_request[i].rd_v.register_value = 'x;
                dispatch_request[i].rd_v.ROB_ID = 'x;
                dispatch_request[i].rd_v.dependency = 'x;
                dispatch_request[i].rd_en = 1'b0;

                // Setup entries going to reservation station
                // ROB Setup
                rs_rob_entry[i].rob.rob_id = 'x;
                rs_rob_entry[i].rob.commit = 'x;
                rs_rob_entry[i].rs_entry.input1_met = 'x;
                rs_rob_entry[i].rs_entry.input2_met = 'x;
                rs_rob_entry[i].rs_entry.rs1_source = 'x;
                rs_rob_entry[i].rs_entry.rs2_source = 'x;
                rs_rob_entry[i].rs_entry.full = 'x;
                rs_rob_entry[i].rob.branch_enable = 'x;
                rs_rob_entry[i].rob.mispredict = '0;
                // RVFI setup
                rs_rob_entry[i].rvfi.valid = 'x; // SOUMIL IS SLOW
                rs_rob_entry[i].rvfi.order = 'x; // SOUMIL IS SLOW // Need to put actual order here
                rs_rob_entry[i].rvfi.inst = 'x;
                rs_rob_entry[i].rvfi.rs1_addr = 'x;
                rs_rob_entry[i].rvfi.rs2_addr = 'x;
                rs_rob_entry[i].rvfi.rs1_rdata = 'x;
                rs_rob_entry[i].rvfi.rs2_rdata = 'x;
                rs_rob_entry[i].rvfi.rd_addr = 'x;
                rs_rob_entry[i].rvfi.rd_wdata = 'x;
                rs_rob_entry[i].rvfi.pc_rdata = 'x;
                rs_rob_entry[i].rvfi.pc_wdata = 'x;
                rs_rob_entry[i].rvfi.mem_addr = 'x;
                // Need to compute rmask/wmask based on type of mem op
                rs_rob_entry[i].rvfi.mem_rmask = 'x;
                rs_rob_entry[i].rvfi.mem_wmask = 'x;
                rs_rob_entry[i].rvfi.mem_rdata = 'x;
                rs_rob_entry[i].rvfi.mem_wdata = 'x;

                //inst setup
                rs_rob_entry[i].inst = 'x;

                //Rat Registers
                rs_rob_entry[i].rat.rs1 = 'x;
                rs_rob_entry[i].rat.rs2 = 'x;
                rs_rob_entry[i].rat.rd = 'x;

                // Set cross tail for load store queue
                rs_rob_entry[i].cross_entry = 'x;
            end
        end
    end
    
endmodule : dispatcher
